`timescale 1ns/1ps

//**************************************************************************
//************** TEST BENCH FOR SIMULATIONS ********************************
//**************************************************************************

`include "parameter.v"

module first_tb;

//---------------------------------------------------------------------------
//----------------  INTERNAL SIGNALS   --------------------------------------
//---------------------------------------------------------------------------

reg clk;
reg reset;
wire [7:0]RED;
wire [7:0]GREEN;
wire [7:0]BLUE;
wire done;

//---------------------------------------------------------------------------
//---------------  DIFFERENT DUT COMPONENTS   -------------------------------
//---------------------------------------------------------------------------

image_read #(.INFILE(`INPUT_FILE))  dutR (.clk(clk),
                                          .reset(reset),
                                          .red(RED),
                                          .green(GREEN),
                                          .blue(BLUE));
					  
image_write #(.INFILE(`OUTPUT_FILE)) dutW(.clk(clk),
                                          .reset(reset),
                                          .in_red(RED),
                                          .in_green(GREEN),
                                          .in_blue(BLUE),
                                          .done(done));
													  
//---------------------------------------------------------------------------
//----------------  TEST VECTORS   ------------------------------------------
//---------------------------------------------------------------------------

always begin
	clk=0;
	#10 clk=1;
	#10;
end

initial begin
	reset=0;
	#30;
	reset=1;
end

endmodule
